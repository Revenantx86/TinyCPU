module pc (
    input  wire       clk,
    input  wire       reset,
    input  wire       jump_en,
    input  wire [7:0] jump_addr,
    output reg  [7:0] pc_out
);



endmodule
