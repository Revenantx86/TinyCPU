module regfile (
    input  wire       clk,
    input  wire       reset,
    input  wire       we,
    input  wire [2:0] r_addr_a,
    input  wire [2:0] r_addr_b,
    input  wire [2:0] w_addr,
    input  wire [7:0] w_data,
    output wire [7:0] r_data_a,
    output wire [7:0] r_data_b
);

  

endmodule